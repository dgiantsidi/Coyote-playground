import lynxTypes::*;
import simTypes::*;

// AXIS Generator
class c_gen;

  // Send to driver (mailbox)
  mailbox gen2drv;

  // Params
  c_struct_t params;

  // Completion
  event done;

  // Stream type
  integer strm_type;

  // Sent data from a previous simulation run
  logic [AXI_DATA_BITS-1:0] tdata [48] = '{
    'hd56d79d3119d7e92e1e27c243ba20d218113bf19d60a7a70fc2b404419cb6cb29089bf780bd801b4bf76ccdce7485267c580baf8f0533e90da549fd529416d11,
    'hcd755690c86a77892be7e229cc369e3bf3550d69931869b2e0a49efa013eb855d5156a2098cf7876eb91ff41f21655143e02ff92c7d5268395acb913e2ff150c,
    'h3fcfad2a06246217a482b6cb1a068f36fff723113d78fd17ccdc36c425c91df4862d3f05e709b9b4cd2a5872da2e051db74bbe11e5d27d0fd89ec5822bff39e8,
    'h30ca3659e2ef7b7af0ca94c3d1f52839175b3bafc5ab272bf0e65775ded50e20cb943fcbab1f6d97e10ed0c438862d8ffa16e760c5c6e9ddfdc63d5c130e123c,
    'hbe411c4a16dcffbea3df5323e07ea1a49cf8795801ee3f8ef8e058dfddc27aa6f9e48665a1f11395e79e48c43f35feb28809b928d6ef454af62431e2baae87b3,
    'hd32ce077d32621b0196d5fafc9024ccdf5ab8292d6ab1b12d6c104798a2a93a9dd7a9f1ec2c2449df2414854eb80eee8f9307bf313febfdc17e94b55f1f9b036,
    'h994d2ef8f79269adfd9b3bcaa72d5b0294c8f92ee1557a87cb91a641f21fd3f6e2c9707f9c45c142db9bb4c1a2a92538fe8c0a08af4be4fe96841f34c0204b46,
    'hbbb66aeec63f503f9d31eeb1d0543802da5b1580f0ececded60f32b8eb6232ecebe43abe2c4501d3fa45054aeef8e2940508b220a9ca30e5f11d2da2fceb582a,
    'he0a238191b909a57c55542ab1538ebaca90090b029c385583765a3d6cb694c6df29009a61b91bd53ddd347d6dd974443b7337bb11bd3e683ed96049714f8c563,
    'hd91ce08afdb6cf7fe21df5d40133ed11d4c01ea89ece79b0186ddedad7e8f37928f6b0d7c34f7c23e8c60e37fcd72b2ff5d7c8d9d51e62b6ef22e5422c1f85a8,
    'hd48875d3c6f39d6b256ca2b8d67ce950ee052e138f8c46d027f923abfe0b8c83d8ee6f5795e05be72e83c5a5eff9a190369dd7799218c7c3cf87c6dee8f4cdc7,
    'h9ee355e3f26d9b34293496eab5b78e5385f90ac2ebb1c591b045fd62e92bc790ec749072bd82d158057190f19ccd4332ff3d351ff2c32c0ae3ba369fcfa74d3f,
    'hd4519350aea1c0f3d2fb7320fe69c184c6ba7cdfce6dc679d0327be5d5e7d1cce7e74414048daca7ae37459ef0d2ab13e6868265cba4cf3e27b08c2ef7149901,
    'hedd5a820fe8609e72307e1043daa467ec2ce290ef0e1c2f0b38acb55b02b61a2bbb7e0d832261e148a1f7b2812a2c76cb529e2178164ad41260be67aa915196c,
    'h00000000000000000000000000000000000000000000000000000000000000000000000000000000c0ffee0123456789deadbeef987654320000000000000000,
    'h00000000000000000000000000000000091d8c99c14209cd861fbc0c2b58ebab6d1fdcd966023ac8f3ca10e3965c695fa363acc18557a68864fc765d1135a126,

    'hc6f28ac03c3cdb3dc525d8563ede34df178e48e9cfb03d9acbf8ab02081455e124ae9254f5759abcf2e589dc0f79f3082b01ab46d6831046952ecc0415349f4c,
    'hef223d90ffa08ed72bd32d509c88b40e0e5952382c2afc78ee4e5691d2998982f1473c9fffa830d82e3a5d7d3bbfc8b6bae3bfd8eea625b9245f2c05b58773e9,
    'h93d7270dfc9ffb63c18550d6095a3f32f5b41b8123e31408f7de1f758a7ce7db06ebdfe21da23cce917c1fbceb3733a61cf73426da3be2a7f900c81f1bb4ac3c,
    'h9b442022eade9e05d8214d06fd47f7b51e48c6f5de1e05161c2b27c11dfc286dcc95d710fa0347efe11ccff4004c9e8811882e06a227dfd1bcdf5878cc493888,
    'hc4ffb9ccdbeb6a1ae64b2d5ace66835bcd7657edf600f20882dcbb3bf69936718e75122cf04a3b52cb89c820d6dd217ce78bdfdc92927fe92b0f6e513797f0b0,
    'hd678bfa89311bb721f5bf820039990a9d2571a871975fad4df36ea5bd2df2effc0baa0eb05e5fd4c2462a64eff77eb88d8bb59e9d950ed0f2e7c88b1c142b562,
    'hd037f163f510fe2ab072070b90eaa8adce03d7abd64f5395e3c349ebbf4d48b5270d267fda22b376ad275ec20eb68ef6af422d1609a096751225e9f318569789,
    'hf3fa1842f5ed164202e12461817840cc21537d381ea56206afd8ff6cf281d775d499990ae43bc25bd19f4160aed1a5c2ca0bc8fbcb9d3d11a0e2961525c7f348,
    'heda2d20930771c39e29f44d9d455cdf51cff49cede952a2c2e88da81994d04141377d26b840a1aad25ccf37483b245b9cb1d57c1aa7ebfd3f38010a08fc58cb1,
    'h240f198cb1b0fa9131f7589bda44e88bc3b7f3da3a32681adba169c6c9ca3101edf906b7f7c4f081fea37ec4f9edc2d9cc396162e3dc7945cb26b23cf40b43de,
    'h8f3e3c58a0cbb7949b02741efec03b073f9c465a3cc368d80c0428c3907e0151e12f713ade3f0b46f2bc1244af1e4508db93f79dadc51d7c9dc1ef0d32112c32,
    'hf2a28ebccc62889a88ea7462a2bc5340ea75a33114961d8db1659705cfe63b7ce1ece569f45456d5f156bc3b9a8f67b532a938243d114030de8f7f41c75d7db3,
    'hba87dde1c4c2b9fc9153541f9dde7c35960f10f493a86519bad8560d1ca961acaeb3a907fdaaef06e3062628f965af48e4f4bc12bd2d670739a33b84354df9bf,
    'hdf762fde15dcb794cb747cd9cfaae51b8da01f2d9312bd80afc7739a8fcb4ac3883c9866b861bf589fe37180fdd4d46a0ad6251af765b442efe7d9438a67c3fc,
    'h00000000000000000000000000000000000000000000000000000000000000000000000000000000c0ffee0123456789deadbeef987654320000000000000001,
    'h00000000000000000000000000000000faddef2d352d0a27c7a860c5df44f31016d30d210d28c97f2a6078573e06609456f6bd570a2ac0d532ea8910fcd44d35,

    'hc3854c22c78db4aafd6bd7a1e9efcf611158149dcd452709cb68de80d9957cc0b635a00db026b0971e86f0e1b7c297dc170f86fc1b422de9bb0e8bdffe730831,
    'hf5dae96e231b5b93e6ce1148e2f4d2ffcb656a18affeeb39ed42c1b792e6166ed7b5f17a36cf260ff5b21148387f53aad848f9bf36739ba81d3405269f369dd0,
    'h9acd41f2c19c61b73cdd0ff714f09f8e1d83ffc986d3ae81dac6c8fa85dca264a41861eeb6096175ba29d69397a75d64e2bb4c9324bd6785cbb2cbd10c71048a,
    'ha614febcaa15404b262f4b1cfc01d4d6a3b6026fb9e1beece744ce2caa1329e6065f3ddcec4d8c2f94bd06a9f9a2d889b3828110faf741fd1556233d0cbc6553,
    'h3d58ed1a96bce45c89b2acdfe6d340abd55465d8dc05db34fe0dce76d685ac6fc1687e84adacd1abe8c57235feceb9699a9d5cafd060fccaedc03a3ac299c51b,
    'h2971c204e1b0d5f6e018cb242d58bf9ce59bff83d30362d6dd08fac6fc190268fc14d6738d15684dd04fc4d5e982fd1bd6ee8c63cff39279abc93d921291d958,
    'h364785dbfd13ea65b19205602269a9d593133b7cc5138240b1a9995f13dddc06ea00aee8ec7e8320f0c01075ff355f76db12d357c52b163fa31dcb90eacb4f72,
    'he8e60d3bbc0f6a001e8ea32f04f698cfe2fb56ed023f3497ea7a463ee3ef746cd91413131c4f6e989a7c5290ff0be280a92b2183ce2ad7a6c97321dcda083093,
    'hc75480a9229103e89e56fc2cc4811c16ad5046ef1bf6812d2b4f563802d36493f540bcf882607aff1931c5deaa7ce25ca6b5c434a8eedb38e9a19eb5cac3da9c,
    'h391c9e161c751f14c5df35dfeb8dd3a5ace618fce4db644a2d73fca1cd8eca70ef8f0617e103d195be19d704df574e8cf54c5e33cc702b0c0f74f36c9037b78b,
    'hcefb0f4ee624ad4f84bdf0ad00f86fba86b15b52fc20f51691bf15b6ce029f94df7351fc889cfb97ef395a0338aebbbe9cada31909221a1fdec94591a6c4963e,
    'hc4ad7054f94dea81e809aafaeb545e6782a4ae36f7fc5da0295d25bed95911edf6a93c4af00d4d5ac1f738a9a94b9c4981532155b94fd8639761d943cd5da001,
    'he28e6247be25f72ae5f80290d8e69490d28219e237dec8318a7cf83009a7cdb7eba3dd482e193a5fce699c5fc8da4c2bcc3aeae8dc63bdd1bb3e3157a2c9911d,
    'h1d3ac56cc573ca2d9edfda5f2f2e93901d75bc99e84046dee2651793ee0c31dc27fe0d94369f9381ccc97bfc2f698abdc042394aabc58412a142b5dff89482d7,
    'h00000000000000000000000000000000000000000000000000000000000000000000000000000000c0ffee0123456789deadbeef987654320000000000000002,
    'h000000000000000000000000000000009d26c5f6b51716a5004e165b2edf953fde93edb4fbeea552e971f13104c2a72d3b67252c978439dd5028630c29c0876a
  };

  //
  // C-tor
  //
  function new(mailbox gen2drv, input integer strm_type, input c_struct_t params);
    this.gen2drv = gen2drv;
    this.params = params;
    this.strm_type = strm_type;
  endfunction

  //
  // Run
  // --------------------------------------------------------------------------
  // This is the function to edit if any custom stimulus is needed.
  // By default it will generate random stimulus n_trs times.
  // --------------------------------------------------------------------------
  //

  task run();
    c_trs trs;

    for(int j = 0; j < 3; j++) begin
      for(int i = 0; i < params.n_trs; i++) begin
        trs = new();
        if(!trs.randomize()) $fatal("ERR:  Generator randomization failed");
        trs.tdata = this.tdata[(params.n_trs * j) + i];
        trs.tlast = i == params.n_trs-1;
        trs.display("Gen");
        gen2drv.put(trs);
      end
    end
    -> done;
  endtask

endclass

// for(int j = 0; j < 3; j++) begin
//   for(int i = 0; i < params.n_trs; i++) begin
//     trs = new();
//     if(!trs.randomize()) $fatal("ERR:  Generator randomization failed");
//     trs.tlast = i == params.n_trs-1;
//     trs.display("Gen");
//     gen2drv.put(trs);
//   end
// end
